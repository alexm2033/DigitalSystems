module challenge_B(output wire Y, input wire A, B ,C );
